module top;
import rv32i_types::*;

reservation_station_itf itf();

testbench tb(.*);

endmodule : top;